`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 03/09/2017 05:34:19 PM
// Design Name:
// Module Name: display
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

(* use_dsp48 = "yes" *) module display #
    (
        // 1280 x 1024 display @ 60 Hz
        parameter PIXELS_HORIZ = 80,
        parameter PIXELS_VERT = 64,
        parameter PIXELS_PER_SQ = PIXELS_VERT * PIXELS_HORIZ,
        parameter statusN = 7,		// bits per status reg
        parameter squareN_row = 16,		// rows
        parameter squareN_col = 16,		// columns
        parameter squareN = squareN_row * squareN_col
    )
    (
        input clk, // 100 mhz clock.
        // assume count from left to right, top to bottom.
        input [squareN - 1:0] statusesIn,
        input [31:0] hund, // score
        input [31:0] ten,  // score
        input [31:0] oned,  // score
        input [11:0] freq,  // freq from 1 to 1024 (this is artificial since we actually only have 512)
        output [3:0] VGA_RED_O,
        output [3:0] VGA_GREEN_O,
        output [3:0] VGA_BLUE_O,
        output VGA_VS,
        output VGA_HS
    );

    wire ready;
    wire[11:0] col_pos;
    wire[11:0] row_pos;
    wire[11:0] colour;

    vga_controller vga_ctrl_inst(
        .pixel_clk(clk),
        .Hsync(VGA_HS),
        .Vsync(VGA_VS),
        .active(ready),
        .Counter_X(col_pos),
        .Counter_Y(row_pos)
    );

    wire [15:0] sq_row_i, sq_col_i;
    
    assign sq_row_i = (row_pos >> 6) << 4;
    assign sq_col_i = (col_pos >> 4) / 5;

    wire square_type;
    assign square_type = statusesIn[sq_row_i + sq_col_i];

    /* blue */
//    localparam[11:0] background[0:(PIXELS_PER_SQ - 1)] = {
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
//    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf 
//    };

    /* duck */
    localparam[11:0] duck[0:(PIXELS_PER_SQ - 1)] = {
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'hfff, 12'h9cf, 12'h9cf, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h9cf, 12'h9cf, 12'h224, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'haaa, 12'h9cf, 12'h000, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h9cf, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'haaa, 12'h664, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h9cf, 12'h444, 12'h000, 12'h9cf, 12'h000, 12'h000, 12'haaa, 12'h9cf, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h9cf, 12'h664, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h9cf, 12'h444, 12'h000, 12'h888, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h000, 12'h000, 12'h9cf, 12'haaa, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'haaa, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h444, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'hccc, 12'h888, 12'h000, 12'h000, 12'h888, 12'h888, 12'h000, 12'h000, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'hfff, 12'h000, 12'h000, 12'h000, 12'h888, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h444, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h668, 12'hccc, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h668, 12'h000, 12'h000, 12'h224, 12'h9cf, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'hfff, 12'h9cf, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h664, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h664, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hcdc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h668, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h444, 12'haaa, 12'hccc, 12'hccc, 12'haaa, 12'h664, 12'h444, 12'h444, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h668, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h668, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h664, 12'h664, 12'hcdc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h668, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h888, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hccc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hfff, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'haaa, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hfff, 12'h000, 12'h000, 12'h000, 12'h000, 12'h224, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h888, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h000, 12'h000, 12'h000, 12'hcdc, 12'h664, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'hcdc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'haaa, 12'h000, 12'h000, 12'hcdc, 12'h9cf, 12'hcdc, 12'h444, 12'h000, 12'h224, 12'h000, 12'h000, 12'h000, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'hcdc, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h444, 12'h9cf, 12'h000, 12'haaa, 12'haaa, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 
    12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf, 12'h9cf
    };
    
    reg [15:0] pic_index = 16'b0;
    reg [15:0] one, two, three, four = 16'b0;
    wire [15:0] delay = 16'b0000000000000011;
    
    always @(posedge clk) begin
        if (ready == 1'b1) begin
            one <= row_pos % PIXELS_VERT;
            two <= col_pos % PIXELS_HORIZ;
            three <= one * PIXELS_HORIZ;
            four <= two + three;
            pic_index <= four + delay;
        end
    end                 
    
//    wire [15:0] fake;
//    assign fake = ((row_pos % PIXELS_VERT) * PIXELS_HORIZ) + col_pos % PIXELS_HORIZ;  

    // Display the score as well
    wire [3:0] hund_red, hund_grn, hund_blu, ten_red, ten_grn, ten_blu, one_red, one_grn, one_blu, lab_red, lab_grn, lab_blu;
    
    disp_score hundreds(
        .pixel_clk(clk),
        .score(hund),
        .index(pic_index),
        .VGA_RED(hund_red),
        .VGA_GREEN(hund_grn),
        .VGA_BLUE(hund_blu)
    );
    
    disp_score tens(
        .pixel_clk(clk),
        .score(ten),
        .index(pic_index),
        .VGA_RED(ten_red),
        .VGA_GREEN(ten_grn),
        .VGA_BLUE(ten_blu)    
    );
    
    disp_score ones(
        .pixel_clk(clk),
        .score(oned),
        .index(pic_index),
        .VGA_RED(one_red),
        .VGA_GREEN(one_grn),
        .VGA_BLUE(one_blu)     
    );
    
    disp_labels label(
        .pixel_clk(clk),
        .index(pic_index),
        .sq_row(sq_row_i),
        .sq_col(sq_col_i),
        .VGA_RED(lab_red),
        .VGA_GREEN(lab_grn),
        .VGA_BLUE(lab_blu)
    );
    
    wire [3:0] active;
    assign active[0] = ready;
    assign active[1] = ready;
    assign active[2] = ready;
    assign active[3] = ready;
    
    assign colour = square_type == 12'b0 ? 12'h9cf : duck[pic_index[12:0]];
    reg [3:0] red, green, blue;

    always @(posedge clk) begin 
        // labels for side of screen
        if (sq_row_i == 16'h0000 || sq_col_i == 16'h0000) begin
            red <= lab_red & active;
            green <= lab_grn & active;
            blue <= lab_blu & active;
        // second bottom row reserved for score, displays up to hundreds digit. sq_row_i is 16 times larger than it should be
        end else if (sq_row_i == 16'h00e0) begin
            if (sq_col_i == 16'h000e) begin           // bottom right for ones digit
                red <= one_red & active;
                green <= one_grn & active;
                blue <= one_blu & active;
            end else if (sq_col_i == 16'h000d) begin  // next is tens digit
                red <= ten_red & active;
                green <= ten_grn & active;
                blue <= ten_blu & active;          
            end else if (sq_col_i == 16'h000c) begin  // last is hundreds digit
                red <= hund_red & active;
                green <= hund_grn & active;
                blue <= hund_blu & active;           
            end else begin                      // all other squares are just blank
                red <= 4'h9 & active;
                green <= 4'hc & active;
                blue <= 4'hf & active;
            end
        // part of bottom row is for frequency display
        end else if (sq_row_i == 16'h00f0) begin
            if ((row_pos > 999) && (col_pos < freq + 2) && (col_pos > freq - 2)) begin
                red <= 4'h0;
                green <= 4'h0;
                blue <= 4'h0;
            end else begin
                red <= 4'h9 & active;
                green <= 4'hc & active;
                blue <= 4'hf & active;
            end
        // otherwise display ducks as usual
        end else begin
            red <= colour[11:8] & active;
            green <= colour[7:4] & active;
            blue <= colour[3:0] & active;
        end
    end
    
    assign VGA_RED_O = red;
    assign VGA_GREEN_O = green;
    assign VGA_BLUE_O = blue;

endmodule