`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/02/2017 04:24:24 PM
// Design Name: 
// Module Name: disp_labels
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module disp_labels # (
        // 64 x 80, minus one. Takes up a square per digit
        parameter PIXELS_PER_SQ = 5119
        )
        (
        input pixel_clk,
        input [15:0] index,
        input [15:0] sq_row,
        input [15:0] sq_col,
        output [3:0] VGA_RED,
        output [3:0] VGA_GREEN,
        output [3:0] VGA_BLUE
        );
        
        localparam[11:0] A[0: PIXELS_PER_SQ ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h864, 12'hfff, 12'hfff, 12'hfff, 12'h467, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hace, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h027, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfa3, 12'h000, 12'h000, 12'h000, 12'h049, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h820, 12'h000, 12'h000, 12'h000, 12'h48c, 12'hffb, 12'h200, 12'h000, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h000, 12'h000, 12'h000, 12'h014, 12'hadf, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h001, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h942, 12'h000, 12'h000, 12'h000, 12'h258, 12'hdff, 12'hfff, 12'heb6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h420, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hffd, 12'h610, 12'h000, 12'h000, 12'h000, 12'h013, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h025, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hb84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h48d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h741, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h520, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h6af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h852, 12'h000, 12'h000, 12'h000, 12'h013, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h961, 12'h000, 12'h000, 12'h000, 12'h139, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h359, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h400, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h521, 12'h000, 12'h000, 12'h000, 12'h025, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc82, 12'h000, 12'h000, 12'h000, 12'h003, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h07c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h100, 12'h000, 12'h000, 12'h000, 12'h038, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h940, 12'h000, 12'h000, 12'h000, 12'h000, 12'h7cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h810, 12'h000, 12'h000, 12'h000, 12'h027, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h700, 12'h000, 12'h000, 12'h000, 12'h002, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb52, 12'h000, 12'h000, 12'h000, 12'h001, 12'h456, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h778, 12'h420, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38e, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h421, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h015, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h741, 12'h000, 12'h000, 12'h000, 12'h124, 12'h799, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h865, 12'h100, 12'h000, 12'h000, 12'h000, 12'h247, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h300, 12'h000, 12'h000, 12'h000, 12'h48c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h630, 12'h000, 12'h000, 12'h000, 12'h012, 12'h8bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h962, 12'h000, 12'h000, 12'h000, 12'h012, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h46a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h400, 12'h000, 12'h000, 12'h000, 12'h138, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h310, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h942, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h710, 12'h000, 12'h000, 12'h000, 12'h015, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h037, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h29e, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h002, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h930, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfa4, 12'h000, 12'h000, 12'h000, 12'h000, 12'h16b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h445, 12'hfff, 12'h544, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h744, 12'hfff, 12'hfff, 12'h544, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam[11:0] sharp[0: PIXELS_PER_SQ ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h844, 12'hfff, 12'h554, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb8, 12'h644, 12'hfff, 12'h554, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h038, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h962, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea4, 12'h000, 12'h000, 12'h000, 12'h27c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h740, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb60, 12'h000, 12'h000, 12'h000, 12'h5ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h630, 12'h000, 12'h000, 12'h001, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h830, 12'h000, 12'h000, 12'h001, 12'h6be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h400, 12'h000, 12'h000, 12'h006, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h710, 12'h000, 12'h000, 12'h003, 12'h9de, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec7, 12'h200, 12'h000, 12'h000, 12'h049, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h026, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb6, 12'h100, 12'h000, 12'h000, 12'h05a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h159, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd83, 12'h000, 12'h000, 12'h000, 12'h39e, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca8, 12'h889, 12'h999, 12'h999, 12'h863, 12'h000, 12'h000, 12'h000, 12'h135, 12'h899, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h999, 12'h630, 12'h000, 12'h000, 12'h000, 12'h369, 12'h999, 12'h998, 12'h89b, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb86, 12'h677, 12'h777, 12'h786, 12'h410, 12'h000, 12'h000, 12'h001, 12'h356, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h764, 12'h000, 12'h000, 12'h000, 12'h013, 12'h777, 12'h777, 12'h776, 12'h689, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h721, 12'h000, 12'h000, 12'h014, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffa, 12'h200, 12'h000, 12'h000, 12'h038, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h035, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb5, 12'h000, 12'h000, 12'h000, 12'h26a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h210, 12'h000, 12'h000, 12'h146, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h59d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea6, 12'h100, 12'h000, 12'h000, 12'h258, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb60, 12'h000, 12'h000, 12'h000, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h100, 12'h000, 12'h000, 12'h46b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h820, 12'h000, 12'h000, 12'h003, 12'h9ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h001, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h014, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h842, 12'h000, 12'h000, 12'h002, 12'h6be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h026, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hccc, 12'hccc, 12'hccc, 12'hdb9, 12'h421, 12'h000, 12'h000, 12'h012, 12'h7ac, 12'hdcc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccd, 12'hda6, 12'h000, 12'h000, 12'h000, 12'h136, 12'habc, 12'hccc, 12'hccc, 12'hdde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h137, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h034, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h544, 12'h334, 12'h444, 12'h321, 12'h000, 12'h000, 12'h000, 12'h012, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h444, 12'h443, 12'h200, 12'h000, 12'h000, 12'h000, 12'h123, 12'h444, 12'h443, 12'h334, 12'h78c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h831, 12'h000, 12'h000, 12'h013, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h000, 12'h000, 12'h000, 12'h38d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h310, 12'h000, 12'h000, 12'h024, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h852, 12'h000, 12'h000, 12'h000, 12'h7cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h210, 12'h000, 12'h000, 12'h035, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h741, 12'h000, 12'h000, 12'h000, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h200, 12'h000, 12'h000, 12'h247, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h620, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea6, 12'h100, 12'h000, 12'h000, 12'h248, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h300, 12'h000, 12'h000, 12'h018, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h100, 12'h000, 12'h000, 12'h46b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec8, 12'h200, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h953, 12'h000, 12'h000, 12'h001, 12'h59d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda5, 12'h000, 12'h000, 12'h000, 12'h06b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h842, 12'h000, 12'h000, 12'h001, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h644, 12'hfff, 12'h544, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hb87, 12'h545, 12'hfff, 12'h667, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] B[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h455, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h544, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h236, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h46a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h17b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h531, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb72, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h600, 12'h000, 12'h000, 12'h000, 12'h029, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd81, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'ha60, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h002, 12'h698, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h875, 12'h100, 12'h000, 12'h000, 12'h000, 12'h012, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h269, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h002, 12'h698, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h889, 12'h630, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hace, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'hddc, 12'h740, 12'h000, 12'h000, 12'h000, 12'h000, 12'h024, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h147, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h842, 12'h000, 12'h000, 12'h000, 12'h014, 12'h9ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h100, 12'h000, 12'h000, 12'h002, 12'h6ac, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h100, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h100, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h410, 12'h000, 12'h000, 12'h000, 12'h013, 12'h9ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h521, 12'h000, 12'h000, 12'h000, 12'h000, 12'h248, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h012, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h024, 12'h9ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h455, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h544, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] C[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haab, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc96, 12'h455, 12'h531, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h246, 12'h554, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h17c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heda, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'ha96, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h542, 12'h000, 12'h000, 12'h001, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h410, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h531, 12'h000, 12'h58c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha31, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'hbbc, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfa5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h941, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h310, 12'h000, 12'h000, 12'h000, 12'h014, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h369, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h530, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdb, 12'h520, 12'h000, 12'h000, 12'h000, 12'h024, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h410, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h300, 12'h000, 12'h000, 12'h000, 12'h135, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb8, 12'h300, 12'h000, 12'h000, 12'h000, 12'h135, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h310, 12'h000, 12'h000, 12'h000, 12'h135, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h410, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdb, 12'h530, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h531, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h852, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha52, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h048, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdbb, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd63, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h258, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h553, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h730, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h100, 12'h000, 12'h000, 12'h369, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h841, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'haa7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h369, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h17c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea6, 12'h445, 12'h543, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h355, 12'h554, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'habc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] D[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h864, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h558, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcde, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h950, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h015, 12'h9bb, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h147, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'h9de, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb9, 12'h642, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hdb7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h27c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h014, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h841, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd96, 12'h200, 12'h000, 12'h000, 12'h000, 12'h248, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h420, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h742, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb64, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb64, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h742, 12'h000, 12'h000, 12'h000, 12'h024, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h420, 12'h000, 12'h000, 12'h000, 12'h135, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h300, 12'h000, 12'h000, 12'h000, 12'h359, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h741, 12'h000, 12'h000, 12'h000, 12'h012, 12'h7bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h115, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hed9, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h129, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heca, 12'h854, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h600, 12'h011, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h259, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h950, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hbbb, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h158, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h864, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h544, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] E[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h468, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h110, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h012, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h222, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h110, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h457, 12'hace, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] F[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdb, 12'h764, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h544, 12'h5ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h963, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h007, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h113, 12'h688, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h887, 12'h79b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h006, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h136, 12'hade, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h752, 12'h000, 12'h000, 12'h000, 12'h237, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h741, 12'h000, 12'h000, 12'h000, 12'h137, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hc98, 12'h545, 12'hfff, 12'hfff, 12'h78c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] G[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc9a, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'ha9b, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha86, 12'h455, 12'h553, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h234, 12'hfff, 12'h456, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h014, 12'h9cd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hca6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h038, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h058, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'h973, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdb, 12'h520, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'h9de, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h950, 12'h000, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h620, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha96, 12'h310, 12'h002, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdc, 12'hbac, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h630, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h026, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h953, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h631, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h310, 12'h000, 12'h000, 12'h000, 12'h258, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda7, 12'h200, 12'h000, 12'h000, 12'h001, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc96, 12'h200, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedb, 12'h977, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h9ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h002, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha63, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h006, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h002, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h962, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda7, 12'h200, 12'h000, 12'h000, 12'h001, 12'h47b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hddd, 12'hb73, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h258, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h420, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h742, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h100, 12'h000, 12'h000, 12'h000, 12'h148, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h310, 12'h000, 12'h000, 12'h000, 12'h000, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h015, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd94, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7ac, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea4, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'h9de, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h200, 12'h000, 12'h000, 12'h000, 12'h002, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h058, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haab, 12'hbba, 12'h731, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedb, 12'h620, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h017, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7bc, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfca, 12'h644, 12'h556, 12'h310, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h344, 12'hfff, 12'h566, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'haac, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] oct_two[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h975, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h845, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h830, 12'h011, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h100, 12'h15b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc73, 12'h111, 12'h110, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h023, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heec, 12'h720, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hc85, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfca, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h247, 12'hacc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'ha85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h027, 12'hbdc, 12'hccc, 12'hccc, 12'hccc, 12'hcd9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h007, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h47c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h211, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h059, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h28e, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda4, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h135, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc83, 12'h000, 12'h237, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc94, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedb, 12'haab, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc70, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h8df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h047, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h920, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h016, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h005, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h530, 12'h000, 12'h000, 12'h000, 12'h011, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hb73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h610, 12'h000, 12'h000, 12'h000, 12'h000, 12'h18d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h000, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda4, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha53, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h28d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h037, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8ce, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h001, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h320, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h521, 12'h000, 12'h000, 12'h000, 12'h000, 12'h258, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h531, 12'h000, 12'h000, 12'h000, 12'h011, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h048, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h420, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h017, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h129, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h930, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h962, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h25a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h16a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h001, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc80, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h100, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb73, 12'h100, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h345, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h431, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb83, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69b, 12'hefe, 12'heee, 12'heee, 12'heee, 12'heee, 12'hefd, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h259, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfe9, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h125, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedc, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hacc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h125, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h720, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha74, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h258, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] oct_three[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h975, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h745, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h830, 12'h011, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h100, 12'h15b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h943, 12'h111, 12'h110, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h011, 12'h102, 12'h68c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heec, 12'h720, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hc85, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfca, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h247, 12'hacc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'ha85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h027, 12'hbdc, 12'hccc, 12'hccc, 12'hccc, 12'hcd9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h039, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h47c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h211, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h059, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda4, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h135, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc83, 12'h000, 12'h258, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc94, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedb, 12'haab, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h000, 12'h007, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc70, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc95, 12'h000, 12'h000, 12'h000, 12'h000, 12'h006, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h006, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h047, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h007, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h920, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h016, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc84, 12'h000, 12'h000, 12'h000, 12'h000, 12'h17c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h530, 12'h000, 12'h000, 12'h000, 12'h011, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h510, 12'h000, 12'h000, 12'h000, 12'h001, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h000, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h542, 12'h000, 12'h000, 12'h000, 12'h000, 12'h037, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha53, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h432, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h147, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h831, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h233, 12'h235, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h431, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'h8bb, 12'haaa, 12'h9ac, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h731, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h233, 12'h48b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea6, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h027, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h822, 12'h110, 12'h000, 12'h000, 12'h000, 12'h000, 12'h015, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h531, 12'h000, 12'h000, 12'h000, 12'h011, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h25a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h420, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h100, 12'h000, 12'h000, 12'h000, 12'h001, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h129, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h420, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h930, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h962, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h642, 12'h000, 12'h000, 12'h000, 12'h000, 12'h239, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h642, 12'h000, 12'h000, 12'h000, 12'h000, 12'h239, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h16a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h530, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc80, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc96, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h789, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h410, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h345, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h431, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha40, 12'h000, 12'h122, 12'h268, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38e, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69b, 12'hefe, 12'heee, 12'heee, 12'heee, 12'heee, 12'hefd, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h259, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha40, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h007, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd82, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h136, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedc, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hacc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h752, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h579, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfec, 12'h852, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h369, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha74, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h258, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he93, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h322, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] oct_four[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h975, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h830, 12'h011, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h100, 12'h15b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h001, 12'h111, 12'h111, 12'h111, 12'h100, 12'h058, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heec, 12'h720, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hc85, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea7, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h247, 12'hacc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'ha85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h520, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h47c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h211, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h963, 12'h000, 12'h000, 12'h000, 12'h017, 12'h882, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda4, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h135, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc95, 12'h100, 12'h000, 12'h000, 12'h000, 12'haff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc94, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h38c, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc70, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h049, 12'heff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he82, 12'h000, 12'h000, 12'h000, 12'h004, 12'hadf, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h047, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h200, 12'h000, 12'h000, 12'h001, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h920, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h016, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h720, 12'h000, 12'h000, 12'h000, 12'h259, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h530, 12'h000, 12'h000, 12'h000, 12'h011, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h024, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb7, 12'h100, 12'h000, 12'h000, 12'h002, 12'h7ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h000, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfea, 12'h520, 12'h000, 12'h000, 12'h000, 12'h15a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha53, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h005, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h410, 12'h000, 12'h000, 12'h000, 12'h18d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha60, 12'h000, 12'h000, 12'h000, 12'h037, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he95, 12'h000, 12'h000, 12'h000, 12'h015, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hff9, 12'h100, 12'h000, 12'h000, 12'h000, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h531, 12'h000, 12'h000, 12'h000, 12'h011, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha30, 12'h000, 12'h000, 12'h000, 12'h36a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc71, 12'h000, 12'h000, 12'h000, 12'h004, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h420, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfe8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h112, 12'h333, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h122, 12'h322, 12'h222, 12'h222, 12'h246, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h129, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h930, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h962, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc7, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h16a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfee, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9de, 12'hfff, 12'hfff, 12'hfee, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc80, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h345, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h431, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69b, 12'hefe, 12'heee, 12'heee, 12'heee, 12'heee, 12'hefd, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h259, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedc, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hacc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb61, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd83, 12'h000, 12'h000, 12'h000, 12'h005, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha74, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h258, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        localparam [11:0] oct_five[0: PIXELS_PER_SQ] = {
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h975, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h69c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h830, 12'h011, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h100, 12'h15b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda7, 12'h300, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h111, 12'h110, 12'h005, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heec, 12'h720, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h26a, 12'heef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h740, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hc85, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h013, 12'h8be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h5bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha73, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h247, 12'hacc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'ha85, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h9ff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h47c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd9, 12'h211, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h8ef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda4, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h135, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h036, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc94, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc70, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h952, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h300, 12'h000, 12'h000, 12'h000, 12'h002, 12'h7be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h510, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h047, 12'hdef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h920, 12'h000, 12'h000, 12'h000, 12'h001, 12'h58b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h300, 12'h000, 12'h000, 12'h000, 12'h016, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'h7bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfda, 12'h530, 12'h000, 12'h000, 12'h000, 12'h011, 12'h9df, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hacf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h5bf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he94, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h853, 12'h000, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h246, 12'h776, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'haef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha53, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h841, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h012, 12'h221, 12'h358, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfed, 12'h840, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h159, 12'hcef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hca8, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h666, 12'h776, 12'h310, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb62, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h37b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfcb, 12'hbbb, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h023, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h359, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h001, 12'h49d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca7, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hd93, 12'h000, 12'h000, 12'h000, 12'h000, 12'h146, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h742, 12'h000, 12'h000, 12'h000, 12'h001, 12'h5ae, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc96, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h7cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hea5, 12'h000, 12'h000, 12'h000, 12'h000, 12'h035, 12'hbdf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfeb, 12'h531, 12'h000, 12'h000, 12'h000, 12'h011, 12'h8cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h741, 12'h000, 12'h000, 12'h000, 12'h000, 12'h38c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h000, 12'h000, 12'h000, 12'h000, 12'h025, 12'hadf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfc9, 12'h420, 12'h000, 12'h000, 12'h000, 12'h014, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h249, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffb, 12'h500, 12'h000, 12'h000, 12'h000, 12'h001, 12'h59c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h129, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h249, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h930, 12'h000, 12'h000, 12'h000, 12'h000, 12'h36a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h962, 12'h000, 12'h000, 12'h000, 12'h000, 12'h4af, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'ha64, 12'h100, 12'h000, 12'h000, 12'h000, 12'h239, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'he92, 12'h000, 12'h000, 12'h000, 12'h000, 12'h004, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec9, 12'h400, 12'h000, 12'h000, 12'h000, 12'h003, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h953, 12'h000, 12'h000, 12'h000, 12'h000, 12'h35a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffc, 12'h400, 12'h000, 12'h000, 12'h000, 12'h000, 12'h16a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h951, 12'h000, 12'h000, 12'h000, 12'h000, 12'h05b, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfdb, 12'h530, 12'h000, 12'h000, 12'h000, 12'h000, 12'h39d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc80, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h6bd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb74, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hc95, 12'h100, 12'h000, 12'h000, 12'h000, 12'h013, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffd, 12'h500, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69d, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'h964, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h3ad, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb8, 12'h789, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heb7, 12'h210, 12'h000, 12'h000, 12'h000, 12'h000, 12'h04a, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hdb6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h001, 12'h345, 12'hbff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfb6, 12'h431, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h15a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha40, 12'h000, 12'h124, 12'h79c, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hb71, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'haff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hda6, 12'h100, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h69b, 12'hefe, 12'heee, 12'heee, 12'heee, 12'heee, 12'hefd, 12'ha64, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h259, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'h940, 12'h000, 12'h000, 12'h000, 12'h000, 12'h003, 12'h9ee, 12'hfee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hffb, 12'h600, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h7cf, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h47a, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h002, 12'h6be, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hedc, 12'h851, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h026, 12'hacc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hec8, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h357, 12'hade, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha50, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h016, 12'hdff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hffe, 12'hca6, 12'h200, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h136, 12'hbef, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'ha74, 12'h223, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h258, 12'hcff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfd8, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h333, 12'h332, 12'h217, 12'heff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
        12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
        };
        
        reg [11:0] colour;
        
        always @ (posedge pixel_clk)
        begin
            case (sq_col[15:0])
                16'h0000:
                begin
                    case (sq_row[15:0])
                        16'h0030: colour <= oct_two[index];
                        16'h0060: colour <= oct_three[index];
                        16'h0090: colour <= oct_four[index];
                        16'h00c0: colour <= oct_five[index];
                        default: colour <= 12'hfff;
                    endcase
                end
                16'h0002: colour <= C[index];
                16'h0003: colour <= sharp[index];
                16'h0004: colour <= D[index];
                16'h0005: colour <= sharp[index];
                16'h0006: colour <= E[index];
                16'h0007: colour <= F[index];
                16'h0008: colour <= sharp[index];
                16'h0009: colour <= G[index];
                16'h000a: colour <= sharp[index];
                16'h000b: colour <= A[index];
                16'h000c: colour <= sharp[index];
                16'h000d: colour <= B[index];
                default: colour <= 12'hfff;
            endcase
        end
        
        assign VGA_RED = colour[11:8];
        assign VGA_GREEN = colour[7:4];
        assign VGA_BLUE = colour[3:0];
        
endmodule