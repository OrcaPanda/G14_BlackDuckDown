`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/23/2017 05:57:32 PM
// Design Name: 
// Module Name: disp_score
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module disp_score # (
        // 64 x 80, minus one. Takes up a square per digit
        parameter PIXELS_PER_SQ = 5119
    )
    (
        input pixel_clk,
        input [31:0] score,
        input [15:0] index,
        output [3:0] VGA_RED,
        output [3:0] VGA_GREEN,
        output [3:0] VGA_BLUE
    );
    
    // The largest-value register corresponds to the top left corner of the screen, while reg0 is the bottom right
    // The score should be in the bottom row at least
    
    // Define the colours for each of the numbers
    localparam[11:0] one_c[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h999, 12'h777, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] two_c[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h777, 12'hfff, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'hfff, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'h999, 12'h999, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h888, 12'h777, 12'h777, 12'h777, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'hfff, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h666, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] three_c[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'hbbb, 12'hccc, 12'hbbb, 12'haaa, 12'h999, 12'h888, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'hddd, 12'hbbb, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'hfff, 12'h444, 12'h333, 12'h333, 12'hfff, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h888, 12'haaa, 12'haaa, 12'h888, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h666, 12'h444, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'hfff, 12'h777, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] four_c[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hddd, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hccc, 12'hddd, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hddd, 12'hccc, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h111, 12'h111, 12'h111, 12'h111, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h222, 12'h111, 12'h222, 12'h222, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h222, 12'h222, 12'h111, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h777, 12'hfff, 12'h666, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h777, 12'h666, 12'h666, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] five[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'h999, 12'h888, 12'h888, 12'h777, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h777, 12'h777, 12'h777, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hbbb, 12'haaa, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hbbb, 12'hccc, 12'hccc, 12'hbbb, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h444, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'hbbb, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] six[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'hfff, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h666, 12'h888, 12'haaa, 12'haaa, 12'haaa, 12'hbbb, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h777, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h888, 12'hbbb, 12'haaa, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h666, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'haaa, 12'h777, 12'hfff, 12'h444, 12'h444, 12'h333, 12'h333, 12'h333, 12'h444, 12'hfff, 12'h666, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] seven[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'haaa, 12'haaa, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'hbbb, 12'haaa, 12'h999, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'haaa, 12'h999, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h999, 12'hbbb, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h222, 12'h222, 12'h222, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h666, 12'h777, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h888, 12'h777, 12'h666, 12'h777, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] eight[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hddd, 12'hddd, 12'hccc, 12'hccc, 12'hddd, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'h444, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h777, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h666, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h888, 12'h666, 12'hfff, 12'h444, 12'h444, 12'h333, 12'h333, 12'h444, 12'h444, 12'hfff, 12'h666, 12'h888, 12'haaa, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] nine[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'heee, 12'heee, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'hfff, 12'h999, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'hddd, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hddd, 12'hccc, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'hbbb, 12'h999, 12'h666, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h444, 12'h222, 12'h333, 12'h444, 12'h333, 12'h444, 12'h444, 12'hfff, 12'h666, 12'h777, 12'h888, 12'h999, 12'hbbb, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff
    };
    
    localparam[11:0] zero[0: PIXELS_PER_SQ ] = {
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h999, 12'h666, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h333, 12'h666, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hccc, 12'haaa, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h444, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h888, 12'hccc, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h777, 12'h333, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'h999, 12'hddd, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h333, 12'haaa, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h777, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h666, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hccc, 12'h888, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h444, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h222, 12'h777, 12'hbbb, 12'heee, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hbbb, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h888, 12'h444, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'hfff, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hbbb, 12'hddd, 12'haaa, 12'h666, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hccc, 12'h666, 12'h222, 12'h111, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h444, 12'hbbb, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hddd, 12'h999, 12'h333, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'hfff, 12'hccc, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'heee, 12'hbbb, 12'h888, 12'hfff, 12'h222, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h000, 12'h111, 12'h222, 12'hfff, 12'h888, 12'hddd, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 
    12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff, 12'hfff 
    };
    
    reg [11:0] colour;
    
    always @ (posedge pixel_clk)
    begin
        case (score[11:8])
            4'h0: colour <= zero[index];
            4'h1: colour <= one_c[index];
            4'h2: colour <= two_c[index];
            4'h3: colour <= three_c[index];
            4'h4: colour <= four_c[index];
            4'h5: colour <= five[index];
            4'h6: colour <= six[index];
            4'h7: colour <= seven[index];
            4'h8: colour <= eight[index];
            4'h9: colour <= nine[index];
            default: colour <= 12'hfff;                       
        endcase      
    end
    
    assign VGA_RED = colour[11:8];
    assign VGA_GREEN = colour[7:4];
    assign VGA_BLUE = colour[3:0];
    
endmodule